module VerilogB
    (
        input b,
        output bb
    );

    assign bb = b;
endmodule : VerilogB