module dti_bypass_register
(
input clk_DR,
input TDI,
input bypass_en,
input captureDR,
output TDO_bypass
);


endmodule