module VerilogA
    (
        input a,
        output aa
    );

    assign aa = a;
endmodule : VerilogA