module b
    (
        input in,
        output out
    );

    assign out = in;
endmodule : b