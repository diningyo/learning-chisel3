module a
    (
        input in,
        output out
    );

    b b (.in(in), .out(out));
endmodule : a